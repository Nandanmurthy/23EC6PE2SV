//------------------------------------------------------------------------------
//File       : dummy_dut.sv
//Author     : Nandan M N/1BM23EC162
//Created    : 2026-02-10
//Module     : dummy_dut
//Project    : SystemVerilog and Verification (23EC6PE2SV)
//Faculty    : Prof. Ajaykumar Devarapalli
//Description: A placeholder dummy DUT for the class-based Packet verification lab.
//------------------------------------------------------------------------------

module dummy_dut;
endmodule
