//------------------------------------------------------------------------------
// File       : alu.sv
// Author     : Nandan M N/1BM23EC162
// Project    : SystemVerilog and Verification (23EC6PE2SV)
// Description: 2-input 8-bit ALU
//------------------------------------------------------------------------------

`timescale 1ns/1ps

package alu_pkg;
  typedef enum bit [1:0] {
    ADD = 0,
    SUB = 1,
    MUL = 2,
    XOR = 3
  } opcode_e;
endpackage

import alu_pkg::*;

module alu (
  input  logic [7:0]  a, b,
  input  opcode_e     op,
  output logic [15:0] result
);

  always_comb begin
    case (op)
      ADD: result = a + b;
      SUB: result = a - b;
      MUL: result = a * b;
      XOR: result = a ^ b;
      default: result = '0;
    endcase
  end

endmodule
